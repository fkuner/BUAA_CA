import RightShifterTypes::*;
import RightShifter::*;

(* synthesize *)
module mkTests (Empty);
   RightShifter logicalShifter <- mkRightShifter;
   RightShifter arithmeticShifter <- mkRightShifter;
   
   // there are many ways to write tests.  Here is a very simple
   // version, just to get you started.
   
   rule test;

      let g = multiplexer1(1, 1, 0);
      if (g != 0) begin
	 $display("result is ", g, " but expected 0");
      end
      else begin
	 $display("correct!");
      end

      let e = multiplexer32(1, 24, 25);
      if (e != 25) begin
    $display("result is ", e, " but expected 0");
      end
      else begin
    $display("correct!");
      end
   
      let c = logicalShifter.shift(LogicalRightShift, 12, 2);
      if (c != 3) begin
	 $display("result is ", c, " but expected 3");
      end
      else begin
	 $display("correct!");
      end

      let b = logicalShifter.shift(LogicalRightShift, 12, 1);
      if (b != 6) begin
	 $display("result is ", b, " but expected 6");
      end
      else begin
	 $display("correct!");
      end

      let a = logicalShifter.shift(LogicalRightShift, 1, 1);
      if (a != 0) begin
	 $display("result is ", a); 
      end
      else begin
	 $display("correct!");
      end
      
      let h = logicalShifter.shift(ArithmeticRightShift, 12, 2);
      if (h != 3) begin
	 $display("result is ", h, " but expected 3");
      end
      else begin
	 $display("correct!");
      end

      let i = logicalShifter.shift(ArithmeticRightShift, -12, 2);
      if (i != -3) begin
	 $display("result is ", i, " but expected -3");
      end
      else begin
	 $display("correct!");
      end

      $finish(0);
   endrule
endmodule
